// *****************************************************************************
// (c) Copyright 2022-2032 , Inc. All rights reserved.
// Module Name  :
// Design Name  :
// Project Name :
// Create Date  : 2022-12-21
// Description  :
//
// *****************************************************************************

// -------------------------------------------------------------------
// Constant Parameter
// -------------------------------------------------------------------

// -------------------------------------------------------------------
// Internal Signals Declarations
// -------------------------------------------------------------------

// -------------------------------------------------------------------
// initial
// -------------------------------------------------------------------
initial begin
  char_x_start = 10'd200;
  char_x_end  = 10'd400;
  char_y_start = 10'd200;
  char_y_end  = 10'd400;
  char_color = 4'd2;
  #100000000
  char_x_start = 10'd100;
  char_x_end  = 10'd150;
  char_y_start = 10'd100;
  char_y_end  = 10'd150;
  char_color = 4'd1;
  #100000000
  $finish;
end

// -------------------------------------------------------------------
// Main Code
// -------------------------------------------------------------------

// -------------------------------------------------------------------
// Assertion Declarations
// -------------------------------------------------------------------
`ifdef SOC_ASSERT_ON

`endif
